module vgactlr();

endmodule
